`define ERR(name) $display("[%4t] Assertion failed: %s", $time, name)
