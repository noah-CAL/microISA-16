//==============================================================================
// SPDX-License-Identifier: AGPL-3.0-or-later
// Copyright (C) 2026 Noah Sedlik
//
// Description:
//
// Notes:
//==============================================================================
import assert_pkg::err;

module cpu_assertions (cpu_if.cpu cpu);
endmodule
