//==============================================================================
// SPDX-License-Identifier: AGPL-3.0-or-later
// Copyright (C) 2026 Noah Sedlik
// 
// Description: 
// Features:
//==============================================================================
module cpu (
  cpu_if.cpu cpu
);
endmodule
