//==============================================================================
// Copyright (C) 2026 Noah Sedlik
// 
// Description: FIFO package defining constants
//==============================================================================
package fifo_pkg;
  parameter DATA_WIDTH = 64;
  parameter FIFO_DEPTH = 512;
endpackage
